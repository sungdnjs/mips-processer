library verilog;
use verilog.vl_types.all;
entity tb_mipscomputer is
end tb_mipscomputer;
